module cpu #(
    parameters
) (
    input logic clock, 
    input logic reset,
    
);
    
endmodule